`include "sample_env.sv"
